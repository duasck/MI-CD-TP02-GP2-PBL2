module main();

	wire x1;
	not x (x1, 1);
	
endmodule
